/* Autogenerate from blif file */

module muxR(
    input   s,
    input   a,
    input   b,
    output  o
);
    assign o = s ? a : b;
endmodule

module bddR(
    input [15:0] in,
    output out
);
    wire w2b088260144, w2b08826015f, w2b088260134, w2b088260185, w2b088260209, w2b08826020b, w2b08826018e, w2b088260130, w2b08826020c, w2b0882601a0, w2b088260179, w2b088260182, w2b0882601a4, w2b08826014c, w2b088260175, w2b088260225, w2b0882601de, w2b08826012e, w2b088260132, w2b088260207, w2b088260163, w2b088260146, w2b08826017a, w2b088260150, w2b0882601ae, w2b088260194, w2b088260184, w2b08826018f, w2b0882601cf, w2b088260210, w2b0882601bf, w2b088260151, w2b08826013f, w2b088260168, w2b0882601fe, w2b088260192, w2b088260178, w2b0882601a7, w2b08826019d, w2b088260133, w2b088260152, w2b0882601b5, w2b088260226, w2b0882601c2, w2b0882601e9, w2b08826020a, w2b0882601be, w2b0882601b3, w2b0882601ef, w2b0882601cc, w2b088260190, w2b088260145, w2b088260167, w2b0882601ed, w2b08826020e, w2b088260136, w2b088260142, w2b08826019e, w2b0882601d4, w2b0882601b4, w2b0882601c3, w2b088260140, w2b0882601e2, w2b0882601fc, w2b088260183, w2b088260161, w2b088260174, w2b088260164, w2b088260176, w2b088260177, w2b0882601ec, w2b0882601fd, w2b088260147, w2b0882601a5, w2b0882601ac, w2b08826011a, w2b0882601f6, w2b08826021a, w2b088260171, w2b08826020f, w2b0882601b6, w2b0882601d2, w2b088260191, w2b08826018a, w2b088260156, w2b0882601e0, w2b088260157, w2b0882601b7, w2b088260160, w2b0882601bd, w2b08826021c, w2b088260208, w2b0882601a3, w2b08826013e, w2b0882601c0, w2b0882601df, w2b08826013d, w2b0882601a6, w2b088260172, w2b08826017b, w2b08826021e, w2b08826012d, w2b0882601c8, w2b0882601cd, w2b0882601d5, w2b0882601f8, w2b0882601d1, w2b0882601e1, w2b0882601a1, w2b0882601f7, w2b088260135, w2b088260218, w2b0882601d3, w2b088260153, w2b08826016e, w2b0882601ce, w2b088260227, w2b0882601e3, w2b088260138, w2b088260193, w2b0882601c1, w2b088260137, w2b088260228, w2b088260141, w2b08826019f, w2b088260155, w2b0882601fa, w2b08826020d, w2b0882601a2, w2b088260131, w2b088260173, w2b088260220, w2b088260219, w2b08826021f, w2b08826021b, w2b0882601ee, w2b0882601e8, w2b088260162, w2b0882601dd, w2b088260195, w2b0882601fb, w2b088260165, w2b088260203, w2b0882601ad, w2b0882601b0, w2b0882601b2, w2b0882601d0, w2b088260166, w2b0882601f9, w2b08826021d, w2b08826012f, w2b08826016d, w2b088260143, w2b0882601b1, w2b088260154;
    muxR m0 (.s(in[15]), .a(w2b08826011a), .b(~w2b08826011a), .o(w2b08826012d));
    muxR m1 (.s(in[14]), .a(w2b08826012d), .b(~w2b08826011a), .o(w2b08826012e));
    muxR m2 (.s(in[13]), .a(w2b08826011a), .b(~w2b08826012e), .o(w2b08826015f));
    muxR m3 (.s(in[12]), .a(w2b08826015f), .b(w2b08826011a), .o(w2b088260218));
    muxR m4 (.s(in[11]), .a(w2b08826011a), .b(w2b088260218), .o(w2b088260219));
    muxR m5 (.s(in[10]), .a(w2b088260219), .b(w2b08826011a), .o(w2b08826021a));
    muxR m6 (.s(in[9]), .a(w2b08826021a), .b(w2b08826011a), .o(w2b08826021b));
    muxR m7 (.s(in[8]), .a(w2b08826021b), .b(w2b08826011a), .o(w2b08826021c));
    muxR m8 (.s(in[7]), .a(w2b08826021c), .b(w2b08826011a), .o(w2b08826021d));
    muxR m9 (.s(in[6]), .a(w2b08826011a), .b(w2b08826021d), .o(w2b08826021e));
    muxR m10 (.s(in[5]), .a(w2b08826021e), .b(w2b08826011a), .o(w2b08826021f));
    muxR m11 (.s(in[4]), .a(w2b08826021f), .b(w2b08826011a), .o(w2b088260220));
    muxR m12 (.s(in[14]), .a(w2b08826011a), .b(~w2b08826012d), .o(w2b088260171));
    muxR m13 (.s(in[13]), .a(w2b08826011a), .b(w2b088260171), .o(w2b088260207));
    muxR m14 (.s(in[12]), .a(w2b08826011a), .b(w2b088260207), .o(w2b088260208));
    muxR m15 (.s(in[11]), .a(w2b088260208), .b(w2b08826011a), .o(w2b088260209));
    muxR m16 (.s(in[10]), .a(w2b08826011a), .b(w2b088260209), .o(w2b08826020a));
    muxR m17 (.s(in[9]), .a(w2b08826011a), .b(w2b08826020a), .o(w2b08826020b));
    muxR m18 (.s(in[8]), .a(w2b08826011a), .b(w2b08826020b), .o(w2b08826020c));
    muxR m19 (.s(in[7]), .a(w2b08826020c), .b(w2b08826011a), .o(w2b08826020d));
    muxR m20 (.s(in[6]), .a(w2b08826020d), .b(w2b08826011a), .o(w2b08826020e));
    muxR m21 (.s(in[5]), .a(w2b08826011a), .b(w2b08826020e), .o(w2b08826020f));
    muxR m22 (.s(in[4]), .a(w2b08826020f), .b(w2b08826011a), .o(w2b088260210));
    muxR m23 (.s(in[3]), .a(w2b088260220), .b(w2b088260210), .o(w2b088260225));
    muxR m24 (.s(in[14]), .a(w2b08826012d), .b(w2b08826011a), .o(w2b08826019d));
    muxR m25 (.s(in[13]), .a(w2b08826019d), .b(w2b08826011a), .o(w2b08826019e));
    muxR m26 (.s(in[12]), .a(w2b08826011a), .b(w2b08826019e), .o(w2b0882601f6));
    muxR m27 (.s(in[11]), .a(w2b08826011a), .b(w2b0882601f6), .o(w2b0882601f7));
    muxR m28 (.s(in[10]), .a(w2b08826011a), .b(w2b0882601f7), .o(w2b0882601f8));
    muxR m29 (.s(in[9]), .a(w2b08826011a), .b(w2b0882601f8), .o(w2b0882601f9));
    muxR m30 (.s(in[8]), .a(w2b0882601f9), .b(w2b08826011a), .o(w2b0882601fa));
    muxR m31 (.s(in[7]), .a(w2b0882601fa), .b(w2b08826011a), .o(w2b0882601fb));
    muxR m32 (.s(in[6]), .a(w2b0882601fb), .b(w2b08826011a), .o(w2b0882601fc));
    muxR m33 (.s(in[5]), .a(w2b08826011a), .b(w2b0882601fc), .o(w2b0882601fd));
    muxR m34 (.s(in[4]), .a(w2b0882601fd), .b(w2b08826011a), .o(w2b0882601fe));
    muxR m35 (.s(in[12]), .a(w2b08826019e), .b(w2b08826011a), .o(w2b08826019f));
    muxR m36 (.s(in[11]), .a(w2b08826019f), .b(w2b08826011a), .o(w2b0882601a0));
    muxR m37 (.s(in[10]), .a(w2b0882601a0), .b(w2b08826011a), .o(w2b0882601a1));
    muxR m38 (.s(in[9]), .a(w2b0882601a1), .b(w2b08826011a), .o(w2b0882601a2));
    muxR m39 (.s(in[8]), .a(w2b08826011a), .b(w2b0882601a2), .o(w2b0882601a3));
    muxR m40 (.s(in[7]), .a(w2b0882601a3), .b(w2b08826011a), .o(w2b0882601ec));
    muxR m41 (.s(in[6]), .a(w2b0882601ec), .b(w2b08826011a), .o(w2b0882601ed));
    muxR m42 (.s(in[5]), .a(w2b08826011a), .b(w2b0882601ed), .o(w2b0882601ee));
    muxR m43 (.s(in[4]), .a(w2b0882601ee), .b(w2b08826011a), .o(w2b0882601ef));
    muxR m44 (.s(in[3]), .a(w2b0882601fe), .b(w2b0882601ef), .o(w2b088260203));
    muxR m45 (.s(in[2]), .a(w2b088260225), .b(w2b088260203), .o(w2b088260226));
    muxR m46 (.s(in[14]), .a(w2b08826011a), .b(w2b08826012d), .o(w2b08826013d));
    muxR m47 (.s(in[13]), .a(w2b08826013d), .b(w2b08826011a), .o(w2b08826013e));
    muxR m48 (.s(in[12]), .a(w2b08826011a), .b(w2b08826013e), .o(w2b08826013f));
    muxR m49 (.s(in[11]), .a(w2b08826011a), .b(w2b08826013f), .o(w2b0882601b0));
    muxR m50 (.s(in[10]), .a(w2b08826011a), .b(w2b0882601b0), .o(w2b0882601dd));
    muxR m51 (.s(in[9]), .a(w2b08826011a), .b(w2b0882601dd), .o(w2b0882601de));
    muxR m52 (.s(in[8]), .a(w2b0882601de), .b(w2b08826011a), .o(w2b0882601df));
    muxR m53 (.s(in[7]), .a(w2b0882601df), .b(w2b08826011a), .o(w2b0882601e0));
    muxR m54 (.s(in[6]), .a(w2b0882601e0), .b(w2b08826011a), .o(w2b0882601e1));
    muxR m55 (.s(in[5]), .a(w2b0882601e1), .b(w2b08826011a), .o(w2b0882601e2));
    muxR m56 (.s(in[4]), .a(w2b08826011a), .b(w2b0882601e2), .o(w2b0882601e3));
    muxR m57 (.s(in[13]), .a(w2b08826011a), .b(w2b08826019d), .o(w2b0882601cc));
    muxR m58 (.s(in[12]), .a(w2b0882601cc), .b(w2b08826011a), .o(w2b0882601cd));
    muxR m59 (.s(in[11]), .a(w2b08826011a), .b(w2b0882601cd), .o(w2b0882601ce));
    muxR m60 (.s(in[10]), .a(w2b0882601ce), .b(w2b08826011a), .o(w2b0882601cf));
    muxR m61 (.s(in[9]), .a(w2b0882601cf), .b(w2b08826011a), .o(w2b0882601d0));
    muxR m62 (.s(in[8]), .a(w2b08826011a), .b(w2b0882601d0), .o(w2b0882601d1));
    muxR m63 (.s(in[7]), .a(w2b08826011a), .b(w2b0882601d1), .o(w2b0882601d2));
    muxR m64 (.s(in[6]), .a(w2b0882601d2), .b(w2b08826011a), .o(w2b0882601d3));
    muxR m65 (.s(in[5]), .a(w2b0882601d3), .b(w2b08826011a), .o(w2b0882601d4));
    muxR m66 (.s(in[4]), .a(w2b0882601d4), .b(w2b08826011a), .o(w2b0882601d5));
    muxR m67 (.s(in[3]), .a(w2b0882601e3), .b(w2b0882601d5), .o(w2b0882601e8));
    muxR m68 (.s(in[12]), .a(w2b08826011a), .b(w2b08826015f), .o(w2b088260160));
    muxR m69 (.s(in[11]), .a(w2b08826011a), .b(w2b088260160), .o(w2b088260161));
    muxR m70 (.s(in[10]), .a(w2b088260161), .b(w2b08826011a), .o(w2b0882601bd));
    muxR m71 (.s(in[9]), .a(w2b0882601bd), .b(w2b08826011a), .o(w2b0882601be));
    muxR m72 (.s(in[8]), .a(w2b08826011a), .b(w2b0882601be), .o(w2b0882601bf));
    muxR m73 (.s(in[7]), .a(w2b0882601bf), .b(w2b08826011a), .o(w2b0882601c0));
    muxR m74 (.s(in[6]), .a(w2b0882601c0), .b(w2b08826011a), .o(w2b0882601c1));
    muxR m75 (.s(in[5]), .a(w2b0882601c1), .b(w2b08826011a), .o(w2b0882601c2));
    muxR m76 (.s(in[4]), .a(w2b0882601c2), .b(w2b08826011a), .o(w2b0882601c3));
    muxR m77 (.s(in[10]), .a(w2b0882601b0), .b(w2b08826011a), .o(w2b0882601b1));
    muxR m78 (.s(in[9]), .a(w2b0882601b1), .b(w2b08826011a), .o(w2b0882601b2));
    muxR m79 (.s(in[8]), .a(w2b08826011a), .b(w2b0882601b2), .o(w2b0882601b3));
    muxR m80 (.s(in[7]), .a(w2b08826011a), .b(w2b0882601b3), .o(w2b0882601b4));
    muxR m81 (.s(in[6]), .a(w2b08826011a), .b(w2b0882601b4), .o(w2b0882601b5));
    muxR m82 (.s(in[5]), .a(w2b08826011a), .b(w2b0882601b5), .o(w2b0882601b6));
    muxR m83 (.s(in[4]), .a(w2b08826011a), .b(w2b0882601b6), .o(w2b0882601b7));
    muxR m84 (.s(in[3]), .a(w2b0882601c3), .b(w2b0882601b7), .o(w2b0882601c8));
    muxR m85 (.s(in[2]), .a(w2b0882601e8), .b(w2b0882601c8), .o(w2b0882601e9));
    muxR m86 (.s(in[1]), .a(w2b088260226), .b(w2b0882601e9), .o(w2b088260227));
    muxR m87 (.s(in[7]), .a(w2b08826011a), .b(w2b0882601a3), .o(w2b0882601a4));
    muxR m88 (.s(in[6]), .a(w2b0882601a4), .b(w2b08826011a), .o(w2b0882601a5));
    muxR m89 (.s(in[5]), .a(w2b08826011a), .b(w2b0882601a5), .o(w2b0882601a6));
    muxR m90 (.s(in[4]), .a(w2b08826011a), .b(w2b0882601a6), .o(w2b0882601a7));
    muxR m91 (.s(in[11]), .a(w2b088260160), .b(w2b08826011a), .o(w2b08826018e));
    muxR m92 (.s(in[10]), .a(w2b08826011a), .b(w2b08826018e), .o(w2b08826018f));
    muxR m93 (.s(in[9]), .a(w2b08826018f), .b(w2b08826011a), .o(w2b088260190));
    muxR m94 (.s(in[8]), .a(w2b08826011a), .b(w2b088260190), .o(w2b088260191));
    muxR m95 (.s(in[7]), .a(w2b088260191), .b(w2b08826011a), .o(w2b088260192));
    muxR m96 (.s(in[6]), .a(w2b088260192), .b(w2b08826011a), .o(w2b088260193));
    muxR m97 (.s(in[5]), .a(w2b08826011a), .b(w2b088260193), .o(w2b088260194));
    muxR m98 (.s(in[4]), .a(w2b08826011a), .b(w2b088260194), .o(w2b088260195));
    muxR m99 (.s(in[3]), .a(w2b0882601a7), .b(w2b088260195), .o(w2b0882601ac));
    muxR m100 (.s(in[13]), .a(w2b08826012e), .b(~w2b08826011a), .o(w2b08826012f));
    muxR m101 (.s(in[12]), .a(w2b08826011a), .b(~w2b08826012f), .o(w2b088260130));
    muxR m102 (.s(in[11]), .a(w2b088260130), .b(w2b08826011a), .o(w2b088260131));
    muxR m103 (.s(in[10]), .a(w2b088260131), .b(w2b08826011a), .o(w2b088260132));
    muxR m104 (.s(in[9]), .a(w2b08826011a), .b(w2b088260132), .o(w2b088260133));
    muxR m105 (.s(in[8]), .a(w2b08826011a), .b(w2b088260133), .o(w2b088260134));
    muxR m106 (.s(in[7]), .a(w2b088260134), .b(w2b08826011a), .o(w2b088260182));
    muxR m107 (.s(in[6]), .a(w2b08826011a), .b(w2b088260182), .o(w2b088260183));
    muxR m108 (.s(in[5]), .a(w2b088260183), .b(w2b08826011a), .o(w2b088260184));
    muxR m109 (.s(in[4]), .a(w2b08826011a), .b(w2b088260184), .o(w2b088260185));
    muxR m110 (.s(in[13]), .a(w2b088260171), .b(w2b08826011a), .o(w2b088260172));
    muxR m111 (.s(in[12]), .a(w2b08826011a), .b(w2b088260172), .o(w2b088260173));
    muxR m112 (.s(in[11]), .a(w2b088260173), .b(w2b08826011a), .o(w2b088260174));
    muxR m113 (.s(in[10]), .a(w2b088260174), .b(w2b08826011a), .o(w2b088260175));
    muxR m114 (.s(in[9]), .a(w2b088260175), .b(w2b08826011a), .o(w2b088260176));
    muxR m115 (.s(in[8]), .a(w2b08826011a), .b(w2b088260176), .o(w2b088260177));
    muxR m116 (.s(in[7]), .a(w2b08826011a), .b(w2b088260177), .o(w2b088260178));
    muxR m117 (.s(in[6]), .a(w2b088260178), .b(w2b08826011a), .o(w2b088260179));
    muxR m118 (.s(in[5]), .a(w2b088260179), .b(w2b08826011a), .o(w2b08826017a));
    muxR m119 (.s(in[4]), .a(w2b08826011a), .b(w2b08826017a), .o(w2b08826017b));
    muxR m120 (.s(in[3]), .a(w2b088260185), .b(w2b08826017b), .o(w2b08826018a));
    muxR m121 (.s(in[2]), .a(w2b0882601ac), .b(w2b08826018a), .o(w2b0882601ad));
    muxR m122 (.s(in[10]), .a(w2b08826011a), .b(w2b088260161), .o(w2b088260162));
    muxR m123 (.s(in[9]), .a(w2b08826011a), .b(w2b088260162), .o(w2b088260163));
    muxR m124 (.s(in[8]), .a(w2b088260163), .b(w2b08826011a), .o(w2b088260164));
    muxR m125 (.s(in[7]), .a(w2b08826011a), .b(w2b088260164), .o(w2b088260165));
    muxR m126 (.s(in[6]), .a(w2b088260165), .b(w2b08826011a), .o(w2b088260166));
    muxR m127 (.s(in[5]), .a(w2b088260166), .b(w2b08826011a), .o(w2b088260167));
    muxR m128 (.s(in[4]), .a(w2b08826011a), .b(w2b088260167), .o(w2b088260168));
    muxR m129 (.s(in[11]), .a(w2b08826011a), .b(w2b088260130), .o(w2b088260150));
    muxR m130 (.s(in[10]), .a(w2b08826011a), .b(w2b088260150), .o(w2b088260151));
    muxR m131 (.s(in[9]), .a(w2b08826011a), .b(w2b088260151), .o(w2b088260152));
    muxR m132 (.s(in[8]), .a(w2b088260152), .b(w2b08826011a), .o(w2b088260153));
    muxR m133 (.s(in[7]), .a(w2b088260153), .b(w2b08826011a), .o(w2b088260154));
    muxR m134 (.s(in[6]), .a(w2b088260154), .b(w2b08826011a), .o(w2b088260155));
    muxR m135 (.s(in[5]), .a(w2b08826011a), .b(w2b088260155), .o(w2b088260156));
    muxR m136 (.s(in[4]), .a(w2b08826011a), .b(w2b088260156), .o(w2b088260157));
    muxR m137 (.s(in[3]), .a(w2b088260168), .b(w2b088260157), .o(w2b08826016d));
    muxR m138 (.s(in[11]), .a(w2b08826013f), .b(w2b08826011a), .o(w2b088260140));
    muxR m139 (.s(in[10]), .a(w2b08826011a), .b(w2b088260140), .o(w2b088260141));
    muxR m140 (.s(in[9]), .a(w2b08826011a), .b(w2b088260141), .o(w2b088260142));
    muxR m141 (.s(in[8]), .a(w2b088260142), .b(w2b08826011a), .o(w2b088260143));
    muxR m142 (.s(in[7]), .a(w2b088260143), .b(w2b08826011a), .o(w2b088260144));
    muxR m143 (.s(in[6]), .a(w2b08826011a), .b(w2b088260144), .o(w2b088260145));
    muxR m144 (.s(in[5]), .a(w2b08826011a), .b(w2b088260145), .o(w2b088260146));
    muxR m145 (.s(in[4]), .a(w2b08826011a), .b(w2b088260146), .o(w2b088260147));
    muxR m146 (.s(in[7]), .a(w2b08826011a), .b(w2b088260134), .o(w2b088260135));
    muxR m147 (.s(in[6]), .a(w2b088260135), .b(w2b08826011a), .o(w2b088260136));
    muxR m148 (.s(in[5]), .a(w2b08826011a), .b(w2b088260136), .o(w2b088260137));
    muxR m149 (.s(in[4]), .a(w2b08826011a), .b(w2b088260137), .o(w2b088260138));
    muxR m150 (.s(in[3]), .a(w2b088260147), .b(w2b088260138), .o(w2b08826014c));
    muxR m151 (.s(in[2]), .a(w2b08826016d), .b(w2b08826014c), .o(w2b08826016e));
    muxR m152 (.s(in[1]), .a(w2b0882601ad), .b(w2b08826016e), .o(w2b0882601ae));
    muxR m153 (.s(in[0]), .a(w2b088260227), .b(w2b0882601ae), .o(w2b088260228));
    assign w2b08826011a = 1;
    assign out = ~w2b088260228;
endmodule