// ethernet_pt.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module ethernet_pt (
		input  wire        clk_clk,                                 //                               clk.clk
		input  wire        reset_reset_n,                           //                             reset.reset_n
		output wire        tse_0_mac_mdio_connection_mdc,           //         tse_0_mac_mdio_connection.mdc
		input  wire        tse_0_mac_mdio_connection_mdio_in,       //                                  .mdio_in
		output wire        tse_0_mac_mdio_connection_mdio_out,      //                                  .mdio_out
		output wire        tse_0_mac_mdio_connection_mdio_oen,      //                                  .mdio_oen
		input  wire        tse_0_mac_misc_connection_ff_tx_crc_fwd, //         tse_0_mac_misc_connection.ff_tx_crc_fwd
		output wire        tse_0_mac_misc_connection_ff_tx_septy,   //                                  .ff_tx_septy
		output wire        tse_0_mac_misc_connection_tx_ff_uflow,   //                                  .tx_ff_uflow
		output wire        tse_0_mac_misc_connection_ff_tx_a_full,  //                                  .ff_tx_a_full
		output wire        tse_0_mac_misc_connection_ff_tx_a_empty, //                                  .ff_tx_a_empty
		output wire [17:0] tse_0_mac_misc_connection_rx_err_stat,   //                                  .rx_err_stat
		output wire [3:0]  tse_0_mac_misc_connection_rx_frm_type,   //                                  .rx_frm_type
		output wire        tse_0_mac_misc_connection_ff_rx_dsav,    //                                  .ff_rx_dsav
		output wire        tse_0_mac_misc_connection_ff_rx_a_full,  //                                  .ff_rx_a_full
		output wire        tse_0_mac_misc_connection_ff_rx_a_empty, //                                  .ff_rx_a_empty
		input  wire [3:0]  tse_0_mac_rgmii_connection_rgmii_in,     //        tse_0_mac_rgmii_connection.rgmii_in
		output wire [3:0]  tse_0_mac_rgmii_connection_rgmii_out,    //                                  .rgmii_out
		input  wire        tse_0_mac_rgmii_connection_rx_control,   //                                  .rx_control
		output wire        tse_0_mac_rgmii_connection_tx_control,   //                                  .tx_control
		input  wire        tse_0_mac_status_connection_set_10,      //       tse_0_mac_status_connection.set_10
		input  wire        tse_0_mac_status_connection_set_1000,    //                                  .set_1000
		output wire        tse_0_mac_status_connection_eth_mode,    //                                  .eth_mode
		output wire        tse_0_mac_status_connection_ena_10,      //                                  .ena_10
		input  wire        tse_0_pcs_mac_rx_clock_connection_clk,   // tse_0_pcs_mac_rx_clock_connection.clk
		input  wire        tse_0_pcs_mac_tx_clock_connection_clk,   // tse_0_pcs_mac_tx_clock_connection.clk
		output wire        tse_1_mac_mdio_connection_mdc,           //         tse_1_mac_mdio_connection.mdc
		input  wire        tse_1_mac_mdio_connection_mdio_in,       //                                  .mdio_in
		output wire        tse_1_mac_mdio_connection_mdio_out,      //                                  .mdio_out
		output wire        tse_1_mac_mdio_connection_mdio_oen,      //                                  .mdio_oen
		input  wire        tse_1_mac_misc_connection_ff_tx_crc_fwd, //         tse_1_mac_misc_connection.ff_tx_crc_fwd
		output wire        tse_1_mac_misc_connection_ff_tx_septy,   //                                  .ff_tx_septy
		output wire        tse_1_mac_misc_connection_tx_ff_uflow,   //                                  .tx_ff_uflow
		output wire        tse_1_mac_misc_connection_ff_tx_a_full,  //                                  .ff_tx_a_full
		output wire        tse_1_mac_misc_connection_ff_tx_a_empty, //                                  .ff_tx_a_empty
		output wire [17:0] tse_1_mac_misc_connection_rx_err_stat,   //                                  .rx_err_stat
		output wire [3:0]  tse_1_mac_misc_connection_rx_frm_type,   //                                  .rx_frm_type
		output wire        tse_1_mac_misc_connection_ff_rx_dsav,    //                                  .ff_rx_dsav
		output wire        tse_1_mac_misc_connection_ff_rx_a_full,  //                                  .ff_rx_a_full
		output wire        tse_1_mac_misc_connection_ff_rx_a_empty, //                                  .ff_rx_a_empty
		input  wire [3:0]  tse_1_mac_rgmii_connection_rgmii_in,     //        tse_1_mac_rgmii_connection.rgmii_in
		output wire [3:0]  tse_1_mac_rgmii_connection_rgmii_out,    //                                  .rgmii_out
		input  wire        tse_1_mac_rgmii_connection_rx_control,   //                                  .rx_control
		output wire        tse_1_mac_rgmii_connection_tx_control,   //                                  .tx_control
		input  wire        tse_1_mac_status_connection_set_10,      //       tse_1_mac_status_connection.set_10
		input  wire        tse_1_mac_status_connection_set_1000,    //                                  .set_1000
		output wire        tse_1_mac_status_connection_eth_mode,    //                                  .eth_mode
		output wire        tse_1_mac_status_connection_ena_10,      //                                  .ena_10
		input  wire        tse_1_pcs_mac_rx_clock_connection_clk,   // tse_1_pcs_mac_rx_clock_connection.clk
		input  wire        tse_1_pcs_mac_tx_clock_connection_clk    // tse_1_pcs_mac_tx_clock_connection.clk
	);

	wire  [31:0] nios2_data_master_readdata;                          // mm_interconnect_0:nios2_data_master_readdata -> nios2:d_readdata
	wire         nios2_data_master_waitrequest;                       // mm_interconnect_0:nios2_data_master_waitrequest -> nios2:d_waitrequest
	wire         nios2_data_master_debugaccess;                       // nios2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_data_master_debugaccess
	wire  [12:0] nios2_data_master_address;                           // nios2:d_address -> mm_interconnect_0:nios2_data_master_address
	wire   [3:0] nios2_data_master_byteenable;                        // nios2:d_byteenable -> mm_interconnect_0:nios2_data_master_byteenable
	wire         nios2_data_master_read;                              // nios2:d_read -> mm_interconnect_0:nios2_data_master_read
	wire         nios2_data_master_write;                             // nios2:d_write -> mm_interconnect_0:nios2_data_master_write
	wire  [31:0] nios2_data_master_writedata;                         // nios2:d_writedata -> mm_interconnect_0:nios2_data_master_writedata
	wire  [31:0] nios2_instruction_master_readdata;                   // mm_interconnect_0:nios2_instruction_master_readdata -> nios2:i_readdata
	wire         nios2_instruction_master_waitrequest;                // mm_interconnect_0:nios2_instruction_master_waitrequest -> nios2:i_waitrequest
	wire  [12:0] nios2_instruction_master_address;                    // nios2:i_address -> mm_interconnect_0:nios2_instruction_master_address
	wire         nios2_instruction_master_read;                       // nios2:i_read -> mm_interconnect_0:nios2_instruction_master_read
	wire  [31:0] mm_interconnect_0_tse_1_control_port_readdata;       // tse_1:reg_data_out -> mm_interconnect_0:tse_1_control_port_readdata
	wire         mm_interconnect_0_tse_1_control_port_waitrequest;    // tse_1:reg_busy -> mm_interconnect_0:tse_1_control_port_waitrequest
	wire   [7:0] mm_interconnect_0_tse_1_control_port_address;        // mm_interconnect_0:tse_1_control_port_address -> tse_1:reg_addr
	wire         mm_interconnect_0_tse_1_control_port_read;           // mm_interconnect_0:tse_1_control_port_read -> tse_1:reg_rd
	wire         mm_interconnect_0_tse_1_control_port_write;          // mm_interconnect_0:tse_1_control_port_write -> tse_1:reg_wr
	wire  [31:0] mm_interconnect_0_tse_1_control_port_writedata;      // mm_interconnect_0:tse_1_control_port_writedata -> tse_1:reg_data_in
	wire  [31:0] mm_interconnect_0_tse_0_control_port_readdata;       // tse_0:reg_data_out -> mm_interconnect_0:tse_0_control_port_readdata
	wire         mm_interconnect_0_tse_0_control_port_waitrequest;    // tse_0:reg_busy -> mm_interconnect_0:tse_0_control_port_waitrequest
	wire   [7:0] mm_interconnect_0_tse_0_control_port_address;        // mm_interconnect_0:tse_0_control_port_address -> tse_0:reg_addr
	wire         mm_interconnect_0_tse_0_control_port_read;           // mm_interconnect_0:tse_0_control_port_read -> tse_0:reg_rd
	wire         mm_interconnect_0_tse_0_control_port_write;          // mm_interconnect_0:tse_0_control_port_write -> tse_0:reg_wr
	wire  [31:0] mm_interconnect_0_tse_0_control_port_writedata;      // mm_interconnect_0:tse_0_control_port_writedata -> tse_0:reg_data_in
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_readdata;    // nios2:debug_mem_slave_readdata -> mm_interconnect_0:nios2_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_debug_mem_slave_waitrequest; // nios2:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_debug_mem_slave_debugaccess; // mm_interconnect_0:nios2_debug_mem_slave_debugaccess -> nios2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_debug_mem_slave_address;     // mm_interconnect_0:nios2_debug_mem_slave_address -> nios2:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_debug_mem_slave_read;        // mm_interconnect_0:nios2_debug_mem_slave_read -> nios2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_debug_mem_slave_byteenable;  // mm_interconnect_0:nios2_debug_mem_slave_byteenable -> nios2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_debug_mem_slave_write;       // mm_interconnect_0:nios2_debug_mem_slave_write -> nios2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_writedata;   // mm_interconnect_0:nios2_debug_mem_slave_writedata -> nios2:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;    // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;      // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [9:0] mm_interconnect_0_onchip_memory2_0_s1_address;       // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;    // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;         // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;     // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;         // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire  [31:0] nios2_irq_irq;                                       // irq_mapper:sender_irq -> nios2:irq
	wire         tse_0_receive_valid;                                 // tse_0:ff_rx_dval -> avalon_st_adapter:in_0_valid
	wire  [31:0] tse_0_receive_data;                                  // tse_0:ff_rx_data -> avalon_st_adapter:in_0_data
	wire         tse_0_receive_ready;                                 // avalon_st_adapter:in_0_ready -> tse_0:ff_rx_rdy
	wire         tse_0_receive_startofpacket;                         // tse_0:ff_rx_sop -> avalon_st_adapter:in_0_startofpacket
	wire         tse_0_receive_endofpacket;                           // tse_0:ff_rx_eop -> avalon_st_adapter:in_0_endofpacket
	wire   [5:0] tse_0_receive_error;                                 // tse_0:rx_err -> avalon_st_adapter:in_0_error
	wire   [1:0] tse_0_receive_empty;                                 // tse_0:ff_rx_mod -> avalon_st_adapter:in_0_empty
	wire         avalon_st_adapter_out_0_valid;                       // avalon_st_adapter:out_0_valid -> tse_1:ff_tx_wren
	wire  [31:0] avalon_st_adapter_out_0_data;                        // avalon_st_adapter:out_0_data -> tse_1:ff_tx_data
	wire         avalon_st_adapter_out_0_ready;                       // tse_1:ff_tx_rdy -> avalon_st_adapter:out_0_ready
	wire         avalon_st_adapter_out_0_startofpacket;               // avalon_st_adapter:out_0_startofpacket -> tse_1:ff_tx_sop
	wire         avalon_st_adapter_out_0_endofpacket;                 // avalon_st_adapter:out_0_endofpacket -> tse_1:ff_tx_eop
	wire         avalon_st_adapter_out_0_error;                       // avalon_st_adapter:out_0_error -> tse_1:ff_tx_err
	wire   [1:0] avalon_st_adapter_out_0_empty;                       // avalon_st_adapter:out_0_empty -> tse_1:ff_tx_mod
	wire         tse_1_receive_valid;                                 // tse_1:ff_rx_dval -> avalon_st_adapter_001:in_0_valid
	wire  [31:0] tse_1_receive_data;                                  // tse_1:ff_rx_data -> avalon_st_adapter_001:in_0_data
	wire         tse_1_receive_ready;                                 // avalon_st_adapter_001:in_0_ready -> tse_1:ff_rx_rdy
	wire         tse_1_receive_startofpacket;                         // tse_1:ff_rx_sop -> avalon_st_adapter_001:in_0_startofpacket
	wire         tse_1_receive_endofpacket;                           // tse_1:ff_rx_eop -> avalon_st_adapter_001:in_0_endofpacket
	wire   [5:0] tse_1_receive_error;                                 // tse_1:rx_err -> avalon_st_adapter_001:in_0_error
	wire   [1:0] tse_1_receive_empty;                                 // tse_1:ff_rx_mod -> avalon_st_adapter_001:in_0_empty
	wire         avalon_st_adapter_001_out_0_valid;                   // avalon_st_adapter_001:out_0_valid -> tse_0:ff_tx_wren
	wire  [31:0] avalon_st_adapter_001_out_0_data;                    // avalon_st_adapter_001:out_0_data -> tse_0:ff_tx_data
	wire         avalon_st_adapter_001_out_0_ready;                   // tse_0:ff_tx_rdy -> avalon_st_adapter_001:out_0_ready
	wire         avalon_st_adapter_001_out_0_startofpacket;           // avalon_st_adapter_001:out_0_startofpacket -> tse_0:ff_tx_sop
	wire         avalon_st_adapter_001_out_0_endofpacket;             // avalon_st_adapter_001:out_0_endofpacket -> tse_0:ff_tx_eop
	wire         avalon_st_adapter_001_out_0_error;                   // avalon_st_adapter_001:out_0_error -> tse_0:ff_tx_err
	wire   [1:0] avalon_st_adapter_001_out_0_empty;                   // avalon_st_adapter_001:out_0_empty -> tse_0:ff_tx_mod
	wire         rst_controller_reset_out_reset;                      // rst_controller:reset_out -> [avalon_st_adapter:in_rst_0_reset, avalon_st_adapter_001:in_rst_0_reset, irq_mapper:reset, mm_interconnect_0:nios2_reset_reset_bridge_in_reset_reset, nios2:reset_n, onchip_memory2_0:reset, rst_translator:in_reset, tse_0:reset, tse_1:reset]
	wire         rst_controller_reset_out_reset_req;                  // rst_controller:reset_req -> [nios2:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]

	ethernet_pt_nios2 nios2 (
		.clk                                 (clk_clk),                                             //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                     //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                           (nios2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_data_master_read),                              //                          .read
		.d_readdata                          (nios2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_data_master_write),                             //                          .write
		.d_writedata                         (nios2_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                    //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                     // custom_instruction_master.readra
	);

	ethernet_pt_onchip_memory2_0 onchip_memory2_0 (
		.clk        (clk_clk),                                          //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	ethernet_pt_tse_0 tse_0 (
		.clk           (clk_clk),                                          // control_port_clock_connection.clk
		.reset         (rst_controller_reset_out_reset),                   //              reset_connection.reset
		.reg_addr      (mm_interconnect_0_tse_0_control_port_address),     //                  control_port.address
		.reg_data_out  (mm_interconnect_0_tse_0_control_port_readdata),    //                              .readdata
		.reg_rd        (mm_interconnect_0_tse_0_control_port_read),        //                              .read
		.reg_data_in   (mm_interconnect_0_tse_0_control_port_writedata),   //                              .writedata
		.reg_wr        (mm_interconnect_0_tse_0_control_port_write),       //                              .write
		.reg_busy      (mm_interconnect_0_tse_0_control_port_waitrequest), //                              .waitrequest
		.tx_clk        (tse_0_pcs_mac_tx_clock_connection_clk),            //   pcs_mac_tx_clock_connection.clk
		.rx_clk        (tse_0_pcs_mac_rx_clock_connection_clk),            //   pcs_mac_rx_clock_connection.clk
		.set_10        (tse_0_mac_status_connection_set_10),               //         mac_status_connection.set_10
		.set_1000      (tse_0_mac_status_connection_set_1000),             //                              .set_1000
		.eth_mode      (tse_0_mac_status_connection_eth_mode),             //                              .eth_mode
		.ena_10        (tse_0_mac_status_connection_ena_10),               //                              .ena_10
		.rgmii_in      (tse_0_mac_rgmii_connection_rgmii_in),              //          mac_rgmii_connection.rgmii_in
		.rgmii_out     (tse_0_mac_rgmii_connection_rgmii_out),             //                              .rgmii_out
		.rx_control    (tse_0_mac_rgmii_connection_rx_control),            //                              .rx_control
		.tx_control    (tse_0_mac_rgmii_connection_tx_control),            //                              .tx_control
		.ff_rx_clk     (clk_clk),                                          //      receive_clock_connection.clk
		.ff_tx_clk     (clk_clk),                                          //     transmit_clock_connection.clk
		.ff_rx_data    (tse_0_receive_data),                               //                       receive.data
		.ff_rx_eop     (tse_0_receive_endofpacket),                        //                              .endofpacket
		.rx_err        (tse_0_receive_error),                              //                              .error
		.ff_rx_mod     (tse_0_receive_empty),                              //                              .empty
		.ff_rx_rdy     (tse_0_receive_ready),                              //                              .ready
		.ff_rx_sop     (tse_0_receive_startofpacket),                      //                              .startofpacket
		.ff_rx_dval    (tse_0_receive_valid),                              //                              .valid
		.ff_tx_data    (avalon_st_adapter_001_out_0_data),                 //                      transmit.data
		.ff_tx_eop     (avalon_st_adapter_001_out_0_endofpacket),          //                              .endofpacket
		.ff_tx_err     (avalon_st_adapter_001_out_0_error),                //                              .error
		.ff_tx_mod     (avalon_st_adapter_001_out_0_empty),                //                              .empty
		.ff_tx_rdy     (avalon_st_adapter_001_out_0_ready),                //                              .ready
		.ff_tx_sop     (avalon_st_adapter_001_out_0_startofpacket),        //                              .startofpacket
		.ff_tx_wren    (avalon_st_adapter_001_out_0_valid),                //                              .valid
		.mdc           (tse_0_mac_mdio_connection_mdc),                    //           mac_mdio_connection.mdc
		.mdio_in       (tse_0_mac_mdio_connection_mdio_in),                //                              .mdio_in
		.mdio_out      (tse_0_mac_mdio_connection_mdio_out),               //                              .mdio_out
		.mdio_oen      (tse_0_mac_mdio_connection_mdio_oen),               //                              .mdio_oen
		.ff_tx_crc_fwd (tse_0_mac_misc_connection_ff_tx_crc_fwd),          //           mac_misc_connection.ff_tx_crc_fwd
		.ff_tx_septy   (tse_0_mac_misc_connection_ff_tx_septy),            //                              .ff_tx_septy
		.tx_ff_uflow   (tse_0_mac_misc_connection_tx_ff_uflow),            //                              .tx_ff_uflow
		.ff_tx_a_full  (tse_0_mac_misc_connection_ff_tx_a_full),           //                              .ff_tx_a_full
		.ff_tx_a_empty (tse_0_mac_misc_connection_ff_tx_a_empty),          //                              .ff_tx_a_empty
		.rx_err_stat   (tse_0_mac_misc_connection_rx_err_stat),            //                              .rx_err_stat
		.rx_frm_type   (tse_0_mac_misc_connection_rx_frm_type),            //                              .rx_frm_type
		.ff_rx_dsav    (tse_0_mac_misc_connection_ff_rx_dsav),             //                              .ff_rx_dsav
		.ff_rx_a_full  (tse_0_mac_misc_connection_ff_rx_a_full),           //                              .ff_rx_a_full
		.ff_rx_a_empty (tse_0_mac_misc_connection_ff_rx_a_empty)           //                              .ff_rx_a_empty
	);

	ethernet_pt_tse_0 tse_1 (
		.clk           (clk_clk),                                          // control_port_clock_connection.clk
		.reset         (rst_controller_reset_out_reset),                   //              reset_connection.reset
		.reg_addr      (mm_interconnect_0_tse_1_control_port_address),     //                  control_port.address
		.reg_data_out  (mm_interconnect_0_tse_1_control_port_readdata),    //                              .readdata
		.reg_rd        (mm_interconnect_0_tse_1_control_port_read),        //                              .read
		.reg_data_in   (mm_interconnect_0_tse_1_control_port_writedata),   //                              .writedata
		.reg_wr        (mm_interconnect_0_tse_1_control_port_write),       //                              .write
		.reg_busy      (mm_interconnect_0_tse_1_control_port_waitrequest), //                              .waitrequest
		.tx_clk        (tse_1_pcs_mac_tx_clock_connection_clk),            //   pcs_mac_tx_clock_connection.clk
		.rx_clk        (tse_1_pcs_mac_rx_clock_connection_clk),            //   pcs_mac_rx_clock_connection.clk
		.set_10        (tse_1_mac_status_connection_set_10),               //         mac_status_connection.set_10
		.set_1000      (tse_1_mac_status_connection_set_1000),             //                              .set_1000
		.eth_mode      (tse_1_mac_status_connection_eth_mode),             //                              .eth_mode
		.ena_10        (tse_1_mac_status_connection_ena_10),               //                              .ena_10
		.rgmii_in      (tse_1_mac_rgmii_connection_rgmii_in),              //          mac_rgmii_connection.rgmii_in
		.rgmii_out     (tse_1_mac_rgmii_connection_rgmii_out),             //                              .rgmii_out
		.rx_control    (tse_1_mac_rgmii_connection_rx_control),            //                              .rx_control
		.tx_control    (tse_1_mac_rgmii_connection_tx_control),            //                              .tx_control
		.ff_rx_clk     (clk_clk),                                          //      receive_clock_connection.clk
		.ff_tx_clk     (clk_clk),                                          //     transmit_clock_connection.clk
		.ff_rx_data    (tse_1_receive_data),                               //                       receive.data
		.ff_rx_eop     (tse_1_receive_endofpacket),                        //                              .endofpacket
		.rx_err        (tse_1_receive_error),                              //                              .error
		.ff_rx_mod     (tse_1_receive_empty),                              //                              .empty
		.ff_rx_rdy     (tse_1_receive_ready),                              //                              .ready
		.ff_rx_sop     (tse_1_receive_startofpacket),                      //                              .startofpacket
		.ff_rx_dval    (tse_1_receive_valid),                              //                              .valid
		.ff_tx_data    (avalon_st_adapter_out_0_data),                     //                      transmit.data
		.ff_tx_eop     (avalon_st_adapter_out_0_endofpacket),              //                              .endofpacket
		.ff_tx_err     (avalon_st_adapter_out_0_error),                    //                              .error
		.ff_tx_mod     (avalon_st_adapter_out_0_empty),                    //                              .empty
		.ff_tx_rdy     (avalon_st_adapter_out_0_ready),                    //                              .ready
		.ff_tx_sop     (avalon_st_adapter_out_0_startofpacket),            //                              .startofpacket
		.ff_tx_wren    (avalon_st_adapter_out_0_valid),                    //                              .valid
		.mdc           (tse_1_mac_mdio_connection_mdc),                    //           mac_mdio_connection.mdc
		.mdio_in       (tse_1_mac_mdio_connection_mdio_in),                //                              .mdio_in
		.mdio_out      (tse_1_mac_mdio_connection_mdio_out),               //                              .mdio_out
		.mdio_oen      (tse_1_mac_mdio_connection_mdio_oen),               //                              .mdio_oen
		.ff_tx_crc_fwd (tse_1_mac_misc_connection_ff_tx_crc_fwd),          //           mac_misc_connection.ff_tx_crc_fwd
		.ff_tx_septy   (tse_1_mac_misc_connection_ff_tx_septy),            //                              .ff_tx_septy
		.tx_ff_uflow   (tse_1_mac_misc_connection_tx_ff_uflow),            //                              .tx_ff_uflow
		.ff_tx_a_full  (tse_1_mac_misc_connection_ff_tx_a_full),           //                              .ff_tx_a_full
		.ff_tx_a_empty (tse_1_mac_misc_connection_ff_tx_a_empty),          //                              .ff_tx_a_empty
		.rx_err_stat   (tse_1_mac_misc_connection_rx_err_stat),            //                              .rx_err_stat
		.rx_frm_type   (tse_1_mac_misc_connection_rx_frm_type),            //                              .rx_frm_type
		.ff_rx_dsav    (tse_1_mac_misc_connection_ff_rx_dsav),             //                              .ff_rx_dsav
		.ff_rx_a_full  (tse_1_mac_misc_connection_ff_rx_a_full),           //                              .ff_rx_a_full
		.ff_rx_a_empty (tse_1_mac_misc_connection_ff_rx_a_empty)           //                              .ff_rx_a_empty
	);

	ethernet_pt_mm_interconnect_0 mm_interconnect_0 (
		.sys_clk_clk_clk                         (clk_clk),                                             //                       sys_clk_clk.clk
		.nios2_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                      // nios2_reset_reset_bridge_in_reset.reset
		.nios2_data_master_address               (nios2_data_master_address),                           //                 nios2_data_master.address
		.nios2_data_master_waitrequest           (nios2_data_master_waitrequest),                       //                                  .waitrequest
		.nios2_data_master_byteenable            (nios2_data_master_byteenable),                        //                                  .byteenable
		.nios2_data_master_read                  (nios2_data_master_read),                              //                                  .read
		.nios2_data_master_readdata              (nios2_data_master_readdata),                          //                                  .readdata
		.nios2_data_master_write                 (nios2_data_master_write),                             //                                  .write
		.nios2_data_master_writedata             (nios2_data_master_writedata),                         //                                  .writedata
		.nios2_data_master_debugaccess           (nios2_data_master_debugaccess),                       //                                  .debugaccess
		.nios2_instruction_master_address        (nios2_instruction_master_address),                    //          nios2_instruction_master.address
		.nios2_instruction_master_waitrequest    (nios2_instruction_master_waitrequest),                //                                  .waitrequest
		.nios2_instruction_master_read           (nios2_instruction_master_read),                       //                                  .read
		.nios2_instruction_master_readdata       (nios2_instruction_master_readdata),                   //                                  .readdata
		.nios2_debug_mem_slave_address           (mm_interconnect_0_nios2_debug_mem_slave_address),     //             nios2_debug_mem_slave.address
		.nios2_debug_mem_slave_write             (mm_interconnect_0_nios2_debug_mem_slave_write),       //                                  .write
		.nios2_debug_mem_slave_read              (mm_interconnect_0_nios2_debug_mem_slave_read),        //                                  .read
		.nios2_debug_mem_slave_readdata          (mm_interconnect_0_nios2_debug_mem_slave_readdata),    //                                  .readdata
		.nios2_debug_mem_slave_writedata         (mm_interconnect_0_nios2_debug_mem_slave_writedata),   //                                  .writedata
		.nios2_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_debug_mem_slave_byteenable),  //                                  .byteenable
		.nios2_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_debug_mem_slave_waitrequest), //                                  .waitrequest
		.nios2_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_debug_mem_slave_debugaccess), //                                  .debugaccess
		.onchip_memory2_0_s1_address             (mm_interconnect_0_onchip_memory2_0_s1_address),       //               onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write               (mm_interconnect_0_onchip_memory2_0_s1_write),         //                                  .write
		.onchip_memory2_0_s1_readdata            (mm_interconnect_0_onchip_memory2_0_s1_readdata),      //                                  .readdata
		.onchip_memory2_0_s1_writedata           (mm_interconnect_0_onchip_memory2_0_s1_writedata),     //                                  .writedata
		.onchip_memory2_0_s1_byteenable          (mm_interconnect_0_onchip_memory2_0_s1_byteenable),    //                                  .byteenable
		.onchip_memory2_0_s1_chipselect          (mm_interconnect_0_onchip_memory2_0_s1_chipselect),    //                                  .chipselect
		.onchip_memory2_0_s1_clken               (mm_interconnect_0_onchip_memory2_0_s1_clken),         //                                  .clken
		.tse_0_control_port_address              (mm_interconnect_0_tse_0_control_port_address),        //                tse_0_control_port.address
		.tse_0_control_port_write                (mm_interconnect_0_tse_0_control_port_write),          //                                  .write
		.tse_0_control_port_read                 (mm_interconnect_0_tse_0_control_port_read),           //                                  .read
		.tse_0_control_port_readdata             (mm_interconnect_0_tse_0_control_port_readdata),       //                                  .readdata
		.tse_0_control_port_writedata            (mm_interconnect_0_tse_0_control_port_writedata),      //                                  .writedata
		.tse_0_control_port_waitrequest          (mm_interconnect_0_tse_0_control_port_waitrequest),    //                                  .waitrequest
		.tse_1_control_port_address              (mm_interconnect_0_tse_1_control_port_address),        //                tse_1_control_port.address
		.tse_1_control_port_write                (mm_interconnect_0_tse_1_control_port_write),          //                                  .write
		.tse_1_control_port_read                 (mm_interconnect_0_tse_1_control_port_read),           //                                  .read
		.tse_1_control_port_readdata             (mm_interconnect_0_tse_1_control_port_readdata),       //                                  .readdata
		.tse_1_control_port_writedata            (mm_interconnect_0_tse_1_control_port_writedata),      //                                  .writedata
		.tse_1_control_port_waitrequest          (mm_interconnect_0_tse_1_control_port_waitrequest)     //                                  .waitrequest
	);

	ethernet_pt_irq_mapper irq_mapper (
		.clk        (clk_clk),                        //       clk.clk
		.reset      (rst_controller_reset_out_reset), // clk_reset.reset
		.sender_irq (nios2_irq_irq)                   //    sender.irq
	);

	ethernet_pt_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (6),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (2),
		.outDataWidth    (32),
		.outChannelWidth (0),
		.outErrorWidth   (1),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (clk_clk),                               // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),        // in_rst_0.reset
		.in_0_data           (tse_0_receive_data),                    //     in_0.data
		.in_0_valid          (tse_0_receive_valid),                   //         .valid
		.in_0_ready          (tse_0_receive_ready),                   //         .ready
		.in_0_startofpacket  (tse_0_receive_startofpacket),           //         .startofpacket
		.in_0_endofpacket    (tse_0_receive_endofpacket),             //         .endofpacket
		.in_0_empty          (tse_0_receive_empty),                   //         .empty
		.in_0_error          (tse_0_receive_error),                   //         .error
		.out_0_data          (avalon_st_adapter_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket),   //         .endofpacket
		.out_0_empty         (avalon_st_adapter_out_0_empty),         //         .empty
		.out_0_error         (avalon_st_adapter_out_0_error)          //         .error
	);

	ethernet_pt_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (6),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (2),
		.outDataWidth    (32),
		.outChannelWidth (0),
		.outErrorWidth   (1),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter_001 (
		.in_clk_0_clk        (clk_clk),                                   // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),            // in_rst_0.reset
		.in_0_data           (tse_1_receive_data),                        //     in_0.data
		.in_0_valid          (tse_1_receive_valid),                       //         .valid
		.in_0_ready          (tse_1_receive_ready),                       //         .ready
		.in_0_startofpacket  (tse_1_receive_startofpacket),               //         .startofpacket
		.in_0_endofpacket    (tse_1_receive_endofpacket),                 //         .endofpacket
		.in_0_empty          (tse_1_receive_empty),                       //         .empty
		.in_0_error          (tse_1_receive_error),                       //         .error
		.out_0_data          (avalon_st_adapter_001_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_001_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_001_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_001_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_001_out_0_endofpacket),   //         .endofpacket
		.out_0_empty         (avalon_st_adapter_001_out_0_empty),         //         .empty
		.out_0_error         (avalon_st_adapter_001_out_0_error)          //         .error
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
